module hawk_controller (
    input 
);
    
endmodule